library verilog;
use verilog.vl_types.all;
entity E3_74153_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end E3_74153_vlg_sample_tst;
