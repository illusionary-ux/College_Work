library verilog;
use verilog.vl_types.all;
entity yufei is
    port(
        y               : out    vl_logic;
        b               : in     vl_logic;
        a               : in     vl_logic
    );
end yufei;
