library verilog;
use verilog.vl_types.all;
entity \2023063114THR\ is
    port(
        Q1              : out    vl_logic;
        CLK             : in     vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic;
        Q4              : out    vl_logic;
        Y1              : out    vl_logic;
        Y2              : out    vl_logic;
        Y3              : out    vl_logic;
        Y4              : out    vl_logic;
        D0              : out    vl_logic;
        D1              : out    vl_logic;
        D2              : out    vl_logic;
        D3              : out    vl_logic;
        D4              : out    vl_logic;
        D5              : out    vl_logic;
        D6              : out    vl_logic;
        H0              : out    vl_logic;
        H1              : out    vl_logic;
        H2              : out    vl_logic;
        H3              : out    vl_logic;
        H4              : out    vl_logic;
        H5              : out    vl_logic;
        H6              : out    vl_logic;
        Q0              : out    vl_logic;
        CLK2            : in     vl_logic;
        Q5              : out    vl_logic;
        Q6              : out    vl_logic;
        Q7              : out    vl_logic
    );
end \2023063114THR\;
