library verilog;
use verilog.vl_types.all;
entity jz24_vlg_vec_tst is
end jz24_vlg_vec_tst;
