library verilog;
use verilog.vl_types.all;
entity THR2023063114 is
    port(
        pin_name1       : out    vl_logic;
        clk             : in     vl_logic;
        pin_name2       : out    vl_logic;
        pin_name3       : out    vl_logic;
        pin_name4       : out    vl_logic
    );
end THR2023063114;
