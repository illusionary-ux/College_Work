library verilog;
use verilog.vl_types.all;
entity E3_74138 is
    port(
        RESULT          : out    vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic
    );
end E3_74138;
