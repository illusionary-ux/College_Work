library verilog;
use verilog.vl_types.all;
entity gate_xor is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        Y               : out    vl_logic
    );
end gate_xor;
