library verilog;
use verilog.vl_types.all;
entity test_74147_vlg_check_tst is
    port(
        AN              : in     vl_logic;
        BN              : in     vl_logic;
        CN              : in     vl_logic;
        DN              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test_74147_vlg_check_tst;
