library verilog;
use verilog.vl_types.all;
entity THR2023063114_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end THR2023063114_vlg_sample_tst;
