library verilog;
use verilog.vl_types.all;
entity THR2023063114_vlg_sample_tst is
    port(
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        a3              : in     vl_logic;
        a4              : in     vl_logic;
        a5              : in     vl_logic;
        a6              : in     vl_logic;
        a7              : in     vl_logic;
        a8              : in     vl_logic;
        a9              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end THR2023063114_vlg_sample_tst;
