library verilog;
use verilog.vl_types.all;
entity mo12_vlg_vec_tst is
end mo12_vlg_vec_tst;
