library verilog;
use verilog.vl_types.all;
entity T_14194 is
    port(
        Q0              : out    vl_logic;
        CC              : in     vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic
    );
end T_14194;
