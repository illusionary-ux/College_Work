library verilog;
use verilog.vl_types.all;
entity test_74147 is
    port(
        CN              : out    vl_logic;
        N1              : in     vl_logic;
        N2              : in     vl_logic;
        N3              : in     vl_logic;
        N6              : in     vl_logic;
        N5              : in     vl_logic;
        N4              : in     vl_logic;
        N9              : in     vl_logic;
        N8              : in     vl_logic;
        N7              : in     vl_logic;
        BN              : out    vl_logic;
        AN              : out    vl_logic;
        DN              : out    vl_logic
    );
end test_74147;
