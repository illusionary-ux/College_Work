library verilog;
use verilog.vl_types.all;
entity gate_xor_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end gate_xor_vlg_check_tst;
