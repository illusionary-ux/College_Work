library verilog;
use verilog.vl_types.all;
entity yufei_vlg_vec_tst is
end yufei_vlg_vec_tst;
