library verilog;
use verilog.vl_types.all;
entity jz24_vlg_check_tst is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        a3              : in     vl_logic;
        a4              : in     vl_logic;
        a5              : in     vl_logic;
        a6              : in     vl_logic;
        a7              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end jz24_vlg_check_tst;
