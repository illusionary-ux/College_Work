library verilog;
use verilog.vl_types.all;
entity test_74138_vlg_check_tst is
    port(
        Y0N             : in     vl_logic;
        Y1N             : in     vl_logic;
        Y2N             : in     vl_logic;
        Y3N             : in     vl_logic;
        Y4N             : in     vl_logic;
        Y5N             : in     vl_logic;
        Y6N             : in     vl_logic;
        Y7N             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test_74138_vlg_check_tst;
