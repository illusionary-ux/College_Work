library verilog;
use verilog.vl_types.all;
entity THR2023063114_vlg_check_tst is
    port(
        LED1            : in     vl_logic;
        LED2            : in     vl_logic;
        LED3            : in     vl_logic;
        LED4            : in     vl_logic;
        OA              : in     vl_logic;
        OB              : in     vl_logic;
        OC              : in     vl_logic;
        OD              : in     vl_logic;
        OE              : in     vl_logic;
        \OF\            : in     vl_logic;
        OG              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end THR2023063114_vlg_check_tst;
