library verilog;
use verilog.vl_types.all;
entity three_vlg_vec_tst is
end three_vlg_vec_tst;
