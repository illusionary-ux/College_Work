library verilog;
use verilog.vl_types.all;
entity THR2023063114_vlg_vec_tst is
end THR2023063114_vlg_vec_tst;
