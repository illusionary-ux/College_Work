library verilog;
use verilog.vl_types.all;
entity f_adder_vlg_vec_tst is
end f_adder_vlg_vec_tst;
