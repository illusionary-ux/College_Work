library verilog;
use verilog.vl_types.all;
entity simu_vlg_vec_tst is
end simu_vlg_vec_tst;
