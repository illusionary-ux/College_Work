library verilog;
use verilog.vl_types.all;
entity cnt4_vlg_vec_tst is
end cnt4_vlg_vec_tst;
