library verilog;
use verilog.vl_types.all;
entity E3_74138_vlg_check_tst is
    port(
        RESULT          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end E3_74138_vlg_check_tst;
