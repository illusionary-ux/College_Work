library verilog;
use verilog.vl_types.all;
entity THR2023063114_vlg_check_tst is
    port(
        SOUT            : in     vl_logic;
        SYNC            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end THR2023063114_vlg_check_tst;
