library verilog;
use verilog.vl_types.all;
entity test_74147_vlg_vec_tst is
end test_74147_vlg_vec_tst;
