library verilog;
use verilog.vl_types.all;
entity test_74138 is
    port(
        Y0N             : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        G1              : in     vl_logic;
        C               : in     vl_logic;
        G2AN            : in     vl_logic;
        G2BN            : in     vl_logic;
        Y1N             : out    vl_logic;
        Y2N             : out    vl_logic;
        Y3N             : out    vl_logic;
        Y4N             : out    vl_logic;
        Y5N             : out    vl_logic;
        Y6N             : out    vl_logic;
        Y7N             : out    vl_logic
    );
end test_74138;
