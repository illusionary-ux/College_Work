library verilog;
use verilog.vl_types.all;
entity jz24 is
    port(
        a0              : out    vl_logic;
        cp              : in     vl_logic;
        ld              : in     vl_logic;
        a1              : out    vl_logic;
        a2              : out    vl_logic;
        a3              : out    vl_logic;
        a4              : out    vl_logic;
        a5              : out    vl_logic;
        a6              : out    vl_logic;
        a7              : out    vl_logic
    );
end jz24;
