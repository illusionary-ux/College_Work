library verilog;
use verilog.vl_types.all;
entity E3_74153_vlg_vec_tst is
end E3_74153_vlg_vec_tst;
