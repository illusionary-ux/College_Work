library verilog;
use verilog.vl_types.all;
entity THR2023063114 is
    port(
        SOUT            : out    vl_logic;
        RES             : in     vl_logic;
        CLK             : in     vl_logic;
        SYNC            : out    vl_logic
    );
end THR2023063114;
