library verilog;
use verilog.vl_types.all;
entity cnt4_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end cnt4_vlg_check_tst;
