library verilog;
use verilog.vl_types.all;
entity T_14194_vlg_vec_tst is
end T_14194_vlg_vec_tst;
