library verilog;
use verilog.vl_types.all;
entity E3_74153 is
    port(
        OUTPUT          : out    vl_logic;
        C               : in     vl_logic;
        B               : in     vl_logic;
        A               : in     vl_logic
    );
end E3_74153;
