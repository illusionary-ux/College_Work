library verilog;
use verilog.vl_types.all;
entity test_74283_vlg_vec_tst is
end test_74283_vlg_vec_tst;
