library verilog;
use verilog.vl_types.all;
entity test_74138_vlg_vec_tst is
end test_74138_vlg_vec_tst;
