library verilog;
use verilog.vl_types.all;
entity T_14194_vlg_sample_tst is
    port(
        CC              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end T_14194_vlg_sample_tst;
