library verilog;
use verilog.vl_types.all;
entity Block2 is
    port(
        Y0N             : out    vl_logic;
        pin_name1       : in     vl_logic;
        Y1N             : out    vl_logic;
        Y2N             : out    vl_logic;
        Y3N             : out    vl_logic;
        Y4N             : out    vl_logic;
        Y5N             : out    vl_logic;
        Y6N             : out    vl_logic;
        Y7N             : out    vl_logic
    );
end Block2;
