library verilog;
use verilog.vl_types.all;
entity THR2023063114 is
    port(
        OB              : out    vl_logic;
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        a3              : in     vl_logic;
        a6              : in     vl_logic;
        a5              : in     vl_logic;
        a4              : in     vl_logic;
        a9              : in     vl_logic;
        a8              : in     vl_logic;
        a7              : in     vl_logic;
        OC              : out    vl_logic;
        OE              : out    vl_logic;
        OD              : out    vl_logic;
        \OF\            : out    vl_logic;
        OG              : out    vl_logic;
        OA              : out    vl_logic;
        LED1            : out    vl_logic;
        LED2            : out    vl_logic;
        LED3            : out    vl_logic;
        LED4            : out    vl_logic
    );
end THR2023063114;
