library verilog;
use verilog.vl_types.all;
entity f_adder_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        sout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end f_adder_vlg_check_tst;
