library verilog;
use verilog.vl_types.all;
entity test_74153_vlg_check_tst is
    port(
        Y1              : in     vl_logic;
        Y2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test_74153_vlg_check_tst;
