library verilog;
use verilog.vl_types.all;
entity gate_xor_vlg_vec_tst is
end gate_xor_vlg_vec_tst;
